* E:\STUDY\3rd Semester\SIMULATION\Ex 2 Fig 3.sch

* Schematics Version 9.2
* Sun Jan 28 11:18:08 2018



** Analysis setup **
.DC  TEMP LIST 
+ 27
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Ex 2 Fig 3.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
