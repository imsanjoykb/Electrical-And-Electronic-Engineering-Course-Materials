* E:\STUDY\3rd Semester\SIMULATION\Ex 4 Fig 1.sch

* Schematics Version 9.2
* Wed Jan 31 16:45:14 2018



** Analysis setup **
.DC LIN V_V2 0 20 0.1 
+ LIN V_V1 -4 0 1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Ex 4 Fig 1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
